module flip

// @[noinit]
pub struct Docs {
	label  string
	topics map[string]string
}
